module power_on_reset_sequence #(
) (
);

endmodule
