// Snthesisable code for IEEE754 SP-floating point arithmatic using DSP48 blocks 
// Single-precision Floating Point[IEEE754] Multipler
module floating_point_multipler (
  input  logic clk,
  input  logic [31:0] a,
  input  logic [31:0] b,
  output logic [31:0] p
);

endmodule
