module xilinx_jtag_controller (
);

endmodule
